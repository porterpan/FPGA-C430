// megafunction wizard: %ALTDQ%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTDQ 

// ============================================================
// File Name: mydq.v
// Megafunction Name(s):
// 			ALTDQ
//
// Simulation Library Files(s):
// 			cycloneive
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Build 178 05/31/2012 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module mydq (
	datain_h,
	datain_l,
	inclock,
	oe,
	outclock,
	dataout_h,
	dataout_l,
	padio)/* synthesis synthesis_clearbox = 1 */;

	input	[7:0]  datain_h;
	input	[7:0]  datain_l;
	input	  inclock;
	input	  oe;
	input	  outclock;
	output	[7:0]  dataout_h;
	output	[7:0]  dataout_l;
	inout	[7:0]  padio;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: DDIOINCLK_INPUT STRING "NEGATED_INCLK"
// Retrieval info: CONSTANT: EXTEND_OE_DISABLE STRING "OFF"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: INVERT_INPUT_CLOCKS STRING "ON"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altdq"
// Retrieval info: CONSTANT: NUMBER_OF_DQ NUMERIC "8"
// Retrieval info: CONSTANT: OE_REG STRING "UNREGISTERED"
// Retrieval info: CONSTANT: POWER_UP_HIGH STRING "OFF"
// Retrieval info: USED_PORT: datain_h 0 0 8 0 INPUT NODEFVAL "datain_h[7..0]"
// Retrieval info: CONNECT: @datain_h 0 0 8 0 datain_h 0 0 8 0
// Retrieval info: USED_PORT: datain_l 0 0 8 0 INPUT NODEFVAL "datain_l[7..0]"
// Retrieval info: CONNECT: @datain_l 0 0 8 0 datain_l 0 0 8 0
// Retrieval info: USED_PORT: dataout_h 0 0 8 0 OUTPUT NODEFVAL "dataout_h[7..0]"
// Retrieval info: CONNECT: dataout_h 0 0 8 0 @dataout_h 0 0 8 0
// Retrieval info: USED_PORT: dataout_l 0 0 8 0 OUTPUT NODEFVAL "dataout_l[7..0]"
// Retrieval info: CONNECT: dataout_l 0 0 8 0 @dataout_l 0 0 8 0
// Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "inclock"
// Retrieval info: CONNECT: @inclock 0 0 0 0 inclock 0 0 0 0
// Retrieval info: USED_PORT: oe 0 0 0 0 INPUT NODEFVAL "oe"
// Retrieval info: CONNECT: @oe 0 0 0 0 oe 0 0 0 0
// Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "outclock"
// Retrieval info: CONNECT: @outclock 0 0 0 0 outclock 0 0 0 0
// Retrieval info: USED_PORT: padio 0 0 8 0 BIDIR NODEFVAL "padio[7..0]"
// Retrieval info: CONNECT: padio 0 0 8 0 @padio 0 0 8 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.cmp TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mydq.ppf TRUE FALSE
// Retrieval info: LIB_FILE: cycloneive
